`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// ECE369 - Computer Architecture
// Laboratory 3 (PreLab)
// Module - InstructionMemory.v
// Description - 32-Bit wide instruction memory.
//
// INPUT:-
// Address: 32-Bit address input port.
//
// OUTPUT:-
// Instruction: 32-Bit output port.
//
// FUNCTIONALITY:-
// Similar to the DataMemory, this module should also be byte-addressed
// (i.e., ignore bits 0 and 1 of 'Address'). All of the instructions will be 
// hard-coded into the instruction memory, so there is no need to write to the 
// InstructionMemory.  The contents of the InstructionMemory is the machine 
// language program to be run on your MIPS processor.
////////////////////////////////////////////////////////////////////////////////


module InstructionMemory(Address, Instruction); 

    input [31:0] Address;        // Input Address 

    output [31:0] Instruction;    // Instruction at memory location Address
		
	reg [31:0] memory[0:299];

	
	


	initial begin
	
	
	//branch test instructions
	/*
	memory[0] = 32'b00110100000001000000000000000000;	//	main:		ori	$a0, $zero, 0
memory[1] = 32'b00001000000000000000000000000100;	//			j	start
memory[2] = 32'b00100000000001001111111111111111;	//			addi	$a0, $zero, -1
memory[3] = 32'b00100000000001001111111111111111;	//			addi	$a0, $zero, -1
memory[4] = 32'b10001100100100000000000000000100;	//	start:		lw	$s0, 4($a0)
memory[5] = 32'b10001100100100000000000000001000;	//			lw	$s0, 8($a0)
memory[6] = 32'b10101100100100000000000000000000;	//			sw	$s0, 0($a0)
memory[7] = 32'b10101100100100000000000000001100;	//			sw	$s0, 12($a0)
memory[8] = 32'b10001100100100010000000000000000;	//			lw	$s1, 0($a0)
memory[9] = 32'b10001100100100100000000000001100;	//			lw	$s2, 12($a0)
memory[10] = 32'b00010010000000000000000000000011;	//			beq	$s0, $zero, branch1
memory[11] = 32'b00000010000000001000100000100000;	//			add	$s1, $s0, $zero
memory[12] = 32'b00010010000100010000000000000001;	//			beq	$s0, $s1, branch1
memory[13] = 32'b00001000000000000000000001000100;	//			j	error
memory[14] = 32'b00000110000000011111111111110111;	//	branch1:	bgez	$s0, start
memory[15] = 32'b00100010000100000000000000000001;	//			addi	$s0, $s0, 1
memory[16] = 32'b00000110000000010000000000000001;	//			bgez	$s0, branch2
memory[17] = 32'b00001000000000000000000001000100;	//			j	error
memory[18] = 32'b00100000000100001111111111111111;	//	branch2:	addi	$s0, $zero, -1
memory[19] = 32'b00000000000100000000100000101010;	//			slt	$at, $zero, $s0
memory[20] = 32'b00010100001000000000000000000100;	//			bne	$at, $zero, branch3
memory[21] = 32'b00100000000100000000000000000001;	//			addi	$s0, $zero, 1
memory[22] = 32'b00000000000100000000100000101010;	//			slt	$at, $zero, $s0
memory[23] = 32'b00010100001000000000000000000001;	//			bne	$at, $zero, branch3
memory[24] = 32'b00001000000000000000000001000100;	//			j	error
memory[25] = 32'b00000110000000000000000000000011;	//	branch3:	bltz	$s0, branch4
memory[26] = 32'b00100000000100001111111111111111;	//			addi	$s0, $zero, -1
memory[27] = 32'b00000110000000000000000000000001;	//			bltz	$s0, branch4
memory[28] = 32'b00001000000000000000000001000100;	//			j	error
memory[29] = 32'b00100000000100011111111111111111;	//	branch4:	addi	$s1, $zero, -1
memory[30] = 32'b00010110000100010000000000000010;	//			bne	$s0, $s1, branch5
memory[31] = 32'b00010110000000000000000000000001;	//			bne	$s0, $zero, branch5
memory[32] = 32'b00001000000000000000000001000100;	//			j	error
memory[33] = 32'b00100000000100000000000010000000;	//	branch5:	addi	$s0, $zero, 128
memory[34] = 32'b10100000100100000000000000000000;	//			sb	$s0, 0($a0)
memory[35] = 32'b10000000100100000000000000000000;	//			lb	$s0, 0($a0)
memory[36] = 32'b00011010000000000000000000000001;	//			blez	$s0, branch6
memory[37] = 32'b00001000000000000000000001000100;	//			j	error
memory[38] = 32'b00100000000100001111111111111111;	//	branch6:	addi	$s0, $zero, -1
memory[39] = 32'b00000000000100001000010000000010;	//			srl	$s0, $s0, 16
memory[40] = 32'b10100100100100000000000000000000;	//			sh	$s0, 0($a0)
memory[41] = 32'b00000000000100001000010000000010;	//			srl	$s0, $s0, 16
memory[42] = 32'b10000100100100000000000000000000;	//			lh	$s0, 0($a0)
memory[43] = 32'b00011010000000000000000000000001;	//			blez	$s0, branch7
memory[44] = 32'b00001000000000000000000001000100;	//			j	error
memory[45] = 32'b00100000000100000000000010000000;	//	branch7:	addi	$s0, $zero, 128
memory[46] = 32'b10100000100100000000000000000000;	//			sb	$s0, 0($a0)
memory[47] = 32'b00000000000100001000010000000010;	//			srl	$s0, $s0, 16
memory[48] = 32'b10010000100100000000000000000000;	//			lbu	$s0, 0($a0)
memory[49] = 32'b00000110000000010000000000000001;	//			bgez	$s0, branch8
memory[50] = 32'b00001000000000000000000001000100;	//			j	error
memory[51] = 32'b00100000000100001111111111111111;	//	branch8:	addi	$s0, $zero, -1
memory[52] = 32'b00000000000100001000010000000010;	//			srl	$s0, $s0, 16
memory[53] = 32'b10100100100100000000000000000000;	//			sh	$s0, 0($a0)
memory[54] = 32'b00000000000100001000010000000010;	//			srl	$s0, $s0, 16
memory[55] = 32'b10010100100100000000000000000000;	//			lhu	$s0, 0($a0)
memory[56] = 32'b00000110000000010000000000000001;	//			bgez	$s0, branch9
memory[57] = 32'b00001000000000000000000001000100;	//			j	error
memory[58] = 32'b00100000000100001111111111111111;	//	branch9:	addi	$s0, $zero, -1
memory[59] = 32'b00111100000100000000000000000001;	//			lui	$s0, 1
memory[60] = 32'b00000110000000010000000000000001;	//			bgez	$s0, branch10
memory[61] = 32'b00001000000000000000000001000100;	//			j	error
memory[62] = 32'b00001000000000000000000001000000;	//	branch10:	j	jump1
memory[63] = 32'b00100010000100001111111111111110;	//			addi	$s0, $s0, -2
memory[64] = 32'b00001100000000000000000001000010;	//	jump1:		jal	jal1
memory[65] = 32'b00001000000000000000000000000100;	//			j	start
memory[66] = 32'b00000011111000000000000000001000;	//	jal1:		jr	$ra
memory[67] = 32'b00001000000000000000000001000100;	//			j	error
memory[68] = 32'b00000000000000000000000000001000;	//	error:		jr	$zero

	*/
	/*R-type test instructions
memory[0] = 32'b00100000000100000000000000000001;	//		addi	$s0, $zero, 1
memory[1] = 32'b00100000000100010000000000000001;	//		addi	$s1, $zero, 1
memory[2] = 32'b00000010000100011000000000100100;	//		and	$s0, $s0, $s1
memory[3] = 32'b00000010000000001000000000100100;	//		and	$s0, $s0, $zero
memory[4] = 32'b00000010001100001000000000100010;	//		sub	$s0, $s1, $s0
memory[5] = 32'b00000010000000001000000000100111;	//		nor	$s0, $s0, $zero
memory[6] = 32'b00000010000000001000000000100111;	//		nor	$s0, $s0, $zero
memory[7] = 32'b00000000000000001000000000100101;	//		or	$s0, $zero, $zero
memory[8] = 32'b00000010001000001000000000100101;	//		or	$s0, $s1, $zero
memory[9] = 32'b00000000000100001000000010000000;	//		sll	$s0, $s0, 2
memory[10] = 32'b00000010001100001000000000000100;	//		sllv	$s0, $s0, $s1
memory[11] = 32'b00000010000000001000000000101010;	//		slt	$s0, $s0, $zero
memory[12] = 32'b00000010000100011000000000101010;	//		slt	$s0, $s0, $s1
memory[13] = 32'b00000000000100011000000001000011;	//		sra	$s0, $s1, 1
memory[14] = 32'b00000000000100011000000000000111;	//		srav	$s0, $s1, $zero
memory[15] = 32'b00000000000100011000000001000010;	//		srl	$s0, $s1, 1
memory[16] = 32'b00000000000100011000000011000000;	//		sll	$s0, $s1, 3
memory[17] = 32'b00000000000100001000000011000010;	//		srl	$s0, $s0, 3
memory[18] = 32'b00000010001100001000000000000100;	//		sllv	$s0, $s0, $s1
memory[19] = 32'b00000010001100001000000000000110;	//		srlv	$s0, $s0, $s1
memory[20] = 32'b00000010000100011000000000100110;	//		xor	$s0, $s0, $s1
memory[21] = 32'b00000010000100011000000000100110;	//		xor	$s0, $s0, $s1
memory[22] = 32'b00100000000100100000000000000100;	//		addi	$s2, $zero, 4
memory[23] = 32'b01110010000100101000000000000010;	//		mul	$s0, $s0, $s2
memory[24] = 32'b00100010000100000000000000000100;	//		addi	$s0, $s0, 4
memory[25] = 32'b00110010000100000000000000000000;	//		andi	$s0, $s0, 0
memory[26] = 32'b00110110000100000000000000000001;	//		ori	$s0, $s0, 1
memory[27] = 32'b00101010000100000000000000000000;	//		slti	$s0, $s0, 0
memory[28] = 32'b00101010000100000000000000000001;	//		slti	$s0, $s0, 1
memory[29] = 32'b00111010000100000000000000000001;	//		xori	$s0, $s0, 1
memory[30] = 32'b00111010000100000000000000000001;	//		xori	$s0, $s0, 1
memory[31] = 32'b00100000000100001111111111111110;	//		addi	$s0, $zero, -2
memory[32] = 32'b00100000000100010000000000000010;	//		addi	$s1, $zero, 2
memory[33] = 32'b00000010001100001001000000101011;	//		sltu	$s2, $s1, $s0
memory[34] = 32'b00101110001100001111111111111110;	//		sltiu	$s0, $s1, -2
memory[35] = 32'b00000010001000001000000000001010;	//		movz	$s0, $s1, $zero
memory[36] = 32'b00000000000100011000000000001011;	//		movn	$s0, $zero, $s1
memory[37] = 32'b00000010001100101000000000100000;	//		add	$s0, $s1, $s2
memory[38] = 32'b00100000000100001111111111111110;	//		addi	$s0, $zero, -2
memory[39] = 32'b00000010001100001000100000100001;	//		addu	$s1, $s1, $s0
memory[40] = 32'b00100000000100011111111111111111;	//		addi	$s1, $zero, -1
memory[41] = 32'b01110010001000001001000000100001;	//		clo	$s2, $s1
memory[42] = 32'b00100000000100010000000000000000;	//		addi	$s1, $zero, 0
memory[43] = 32'b01110010001000001001000000100000;	//		clz	$s2, $s1
*/

//GOL
	

	memory[0] = 32'b00000000000000000000000000000000;	//	main:			nop
memory[1] = 32'b00110100000001000000000000000000;	//				ori	$a0, $zero, 0
memory[2] = 32'b00110100000001010000000000010100;	//				ori	$a1, $zero, 20
memory[3] = 32'b00110100000000100000000000000000;	//				ori	$v0, $zero, 0
memory[4] = 32'b00110100000000110000000000000000;	//				ori	$v1, $zero, 0
memory[5] = 32'b00001100000000000000000000000111;	//				jal	gol
memory[6] = 32'b00001000000000000000000000000110;	//	exit:			j	exit
memory[7] = 32'b00110100000010001111111111001110;	//	gol:			ori	$t0, $zero, -50
memory[8] = 32'b00000000000010000100000010000000;	//				sll	$t0, $t0, 2
memory[9] = 32'b00000011101010001110100000100001;	//				addu	$sp, $sp, $t0
memory[10] = 32'b00000011101000000011000000100000;	//				add	$a2, $sp, $zero
memory[11] = 32'b10001100100100000000000000000000;	//				lw	$s0, 0($a0)
memory[12] = 32'b10001100100100010000000000000100;	//				lw	$s1, 4($a0)
memory[13] = 32'b10001100100100100000000000001000;	//				lw	$s2, 8($a0)
memory[14] = 32'b00110100000100110000000000000000;	//				ori	$s3, $zero, 0
memory[15] = 32'b00110100000010000000000000000000;	//				ori	$t0, $zero, 0
memory[16] = 32'b00110100000010100000000000101000;	//				ori	$t2, $zero, 40
memory[17] = 32'b00000000000010000100100010000000;	//	inilizeupdate:		sll	$t1, $t0, 2
memory[18] = 32'b00000001001001100100100000100001;	//				addu	$t1, $t1, $a2
memory[19] = 32'b10101101001000000000000000000000;	//				sw	$zero, 0($t1)
memory[20] = 32'b00100101000010000000000000000001;	//				addiu	$t0, $t0, 1
memory[21] = 32'b00010101000010101111111111111011;	//				bne	$t0, $t2, inilizeupdate
memory[22] = 32'b00000010001000000100000000100000;	//				add	$t0, $s1, $zero
memory[23] = 32'b00100110011100110000000000000001;	//	countcolumns:		addiu	$s3, $s3, 1
memory[24] = 32'b00100101000010001111111111100000;	//				addiu	$t0, $t0, -32
memory[25] = 32'b00010101000000001111111111111101;	//				bne	$t0, $zero, countcolumns
memory[26] = 32'b00110100000101000000000000000000;	//	generation:		ori	$s4, $zero, 0
memory[27] = 32'b00110100000101010000000000000000;	//				ori	$s5, $zero, 0
memory[28] = 32'b00110100000101100000000000000000;	//				ori	$s6, $zero, 0
memory[29] = 32'b00110100000101110000000000000000;	//				ori	$s7, $zero, 0
memory[30] = 32'b01110010100100110100000000000010;	//	getword:		mul	$t0, $s4, $s3
memory[31] = 32'b00000001000101100100000000100001;	//				addu	$t0, $t0, $s6
memory[32] = 32'b00000000000010000100000010000000;	//				sll	$t0, $t0, 2
memory[33] = 32'b00000001000001010100000000100001;	//				addu	$t0, $t0, $a1
memory[34] = 32'b10001101000110010000000000000000;	//				lw	$t9, 0($t0)
memory[35] = 32'b00010110100000000000000000000111;	//	getregisters:		bne	$s4, $zero, nottop
memory[36] = 32'b00100110000010001111111111111111;	//				addiu	$t0, $s0, -1
memory[37] = 32'b01110001000100110100000000000010;	//				mul	$t0, $t0, $s3
memory[38] = 32'b00000001000101100100000000100001;	//				addu	$t0, $t0, $s6
memory[39] = 32'b00000000000010000100000010000000;	//				sll	$t0, $t0, 2
memory[40] = 32'b00000001000001010100000000100001;	//				addu	$t0, $t0, $a1
memory[41] = 32'b10001101000110000000000000000000;	//				lw	$t8, 0($t0)
memory[42] = 32'b00001000000000000000000000110111;	//				j	notbottom
memory[43] = 32'b00100110100010001111111111111111;	//	nottop:			addiu	$t0, $s4, -1
memory[44] = 32'b01110001000100110100000000000010;	//				mul	$t0, $t0, $s3
memory[45] = 32'b00000001000101100100000000100001;	//				addu	$t0, $t0, $s6
memory[46] = 32'b00000000000010000100000010000000;	//				sll	$t0, $t0, 2
memory[47] = 32'b00000001000001010100000000100001;	//				addu	$t0, $t0, $a1
memory[48] = 32'b10001101000110000000000000000000;	//				lw	$t8, 0($t0)
memory[49] = 32'b00100110000010001111111111111111;	//	ifbottom:		addiu	$t0, $s0, -1
memory[50] = 32'b00010101000101000000000000000100;	//				bne	$t0, $s4, notbottom
memory[51] = 32'b00000000000101100100000010000000;	//				sll	$t0, $s6, 2
memory[52] = 32'b00000001000001010100000000100001;	//				addu	$t0, $t0, $a1
memory[53] = 32'b10001101000011110000000000000000;	//				lw	$t7, 0($t0)
memory[54] = 32'b00001000000000000000000000111101;	//				j	ifoleft
memory[55] = 32'b00100110100010000000000000000001;	//	notbottom:		addiu	$t0, $s4, 1
memory[56] = 32'b01110001000100110100000000000010;	//				mul	$t0, $t0, $s3
memory[57] = 32'b00000001000101100100000000100001;	//				addu	$t0, $t0, $s6
memory[58] = 32'b00000000000010000100000010000000;	//				sll	$t0, $t0, 2
memory[59] = 32'b00000001000001010100000000100001;	//				addu	$t0, $t0, $a1
memory[60] = 32'b10001101000011110000000000000000;	//				lw	$t7, 0($t0)
memory[61] = 32'b00010110101000000000000000010100;	//	ifoleft:		bne	$s5, $zero, iforight
memory[62] = 32'b00010110110000000000000000010011;	//				bne	$s6, $zero, iforight
memory[63] = 32'b00100110011010111111111111111111;	//				addiu	$t3, $s3, -1
memory[64] = 32'b01110010100100110100000000000010;	//				mul	$t0, $s4, $s3
memory[65] = 32'b00000001000010110100000000100001;	//				addu	$t0, $t0, $t3
memory[66] = 32'b00010110100000000000000000000100;	//				bne	$s4, $zero, oleftnottop
memory[67] = 32'b00100110000010011111111111111111;	//				addiu	$t1, $s0, -1
memory[68] = 32'b01110001001100110100100000000010;	//				mul	$t1, $t1, $s3
memory[69] = 32'b00000001001010110100100000100001;	//				addu	$t1, $t1, $t3
memory[70] = 32'b00001000000000000000000001001110;	//				j	oleftnotbottom
memory[71] = 32'b00100110100010011111111111111111;	//	oleftnottop:		addiu	$t1, $s4, -1
memory[72] = 32'b01110001001100110100100000000010;	//				mul	$t1, $t1, $s3
memory[73] = 32'b00000001001010110100100000100001;	//				addu	$t1, $t1, $t3
memory[74] = 32'b00100110000010101111111111111111;	//	ifoleftbottom:		addiu	$t2, $s0, -1
memory[75] = 32'b00010101010101000000000000000010;	//				bne	$t2, $s4, oleftnotbottom
memory[76] = 32'b00000001011000000101000000100000;	//				add	$t2, $t3, $zero
memory[77] = 32'b00001000000000000000000010001010;	//				j	end
memory[78] = 32'b00100110100010100000000000000001;	//	oleftnotbottom:		addiu	$t2, $s4, 1
memory[79] = 32'b01110001010100110101000000000010;	//				mul	$t2, $t2, $s3
memory[80] = 32'b00000001010010110101000000100001;	//				addu	$t2, $t2, $t3
memory[81] = 32'b00001000000000000000000010001010;	//				j	end
memory[82] = 32'b00110100000010000000000000011111;	//	iforight:		ori	$t0, $zero, 31
memory[83] = 32'b00100110011010011111111111111111;	//				addiu	$t1, $s3, -1
memory[84] = 32'b00010110101010000000000000001111;	//				bne	$s5, $t0, ifileft
memory[85] = 32'b00010110110010010000000000001110;	//				bne	$s6, $t1, ifileft
memory[86] = 32'b01110010100100110100000000000010;	//				mul	$t0, $s4, $s3
memory[87] = 32'b00010110100000000000000000000011;	//				bne	$s4, $zero, orightnottop
memory[88] = 32'b00100110000010011111111111111111;	//				addiu	$t1, $s0, -1
memory[89] = 32'b01110001001100110100100000000010;	//				mul	$t1, $t1, $s3
memory[90] = 32'b00001000000000000000000001100001;	//				j	orightnotbottom
memory[91] = 32'b00100110100010011111111111111111;	//	orightnottop:		addiu	$t1, $s4, -1
memory[92] = 32'b01110001001100110100100000000010;	//				mul	$t1, $t1, $s3
memory[93] = 32'b00100110000010101111111111111111;	//	iforightbottom:		addiu	$t2, $s0, -1
memory[94] = 32'b00010101010101000000000000000010;	//				bne	$t2, $s4, orightnotbottom
memory[95] = 32'b00110100000010100000000000000000;	//				ori	$t2, $zero, 0
memory[96] = 32'b00001000000000000000000010001010;	//				j	end
memory[97] = 32'b00100110100010100000000000000001;	//	orightnotbottom:	addiu	$t2, $s4, 1
memory[98] = 32'b01110001010100110101000000000010;	//				mul	$t2, $t2, $s3
memory[99] = 32'b00001000000000000000000010001010;	//				j	end
memory[100] = 32'b00010110101000000000000000010011;	//	ifileft:		bne	$s5, $zero, ifiright
memory[101] = 32'b00100110110010111111111111111111;	//				addiu	$t3, $s6, -1
memory[102] = 32'b01110010100100110100000000000010;	//				mul	$t0, $s4, $s3
memory[103] = 32'b00000001000010110100000000100001;	//				addu	$t0, $t0, $t3
memory[104] = 32'b00010110100000000000000000000100;	//				bne	$s4, $zero, ileftnottop
memory[105] = 32'b00100110000010011111111111111111;	//				addiu	$t1, $s0, -1
memory[106] = 32'b01110001001100110100100000000010;	//				mul	$t1, $t1, $s3
memory[107] = 32'b00000001001010110100100000100001;	//				addu	$t1, $t1, $t3
memory[108] = 32'b00001000000000000000000001110100;	//				j	ileftnotbottom
memory[109] = 32'b00100110100010011111111111111111;	//	ileftnottop:		addiu	$t1, $s4, -1
memory[110] = 32'b01110001001100110100100000000010;	//				mul	$t1, $t1, $s3
memory[111] = 32'b00000001001010110100100000100001;	//				addu	$t1, $t1, $t3
memory[112] = 32'b00100110000010101111111111111111;	//	ifileftbottom:		addiu	$t2, $s0, -1
memory[113] = 32'b00010101010101000000000000000010;	//				bne	$t2, $s4, ileftnotbottom
memory[114] = 32'b00000001011000000101000000100000;	//				add	$t2, $t3, $zero
memory[115] = 32'b00001000000000000000000010001010;	//				j	end
memory[116] = 32'b00100110100010100000000000000001;	//	ileftnotbottom:		addiu	$t2, $s4, 1
memory[117] = 32'b01110001010100110101000000000010;	//				mul	$t2, $t2, $s3
memory[118] = 32'b00000001010010110101000000100001;	//				addu	$t2, $t2, $t3
memory[119] = 32'b00001000000000000000000010001010;	//				j	end
memory[120] = 32'b00100110110010110000000000000001;	//	ifiright:		addiu	$t3, $s6, 1
memory[121] = 32'b01110010100100110100000000000010;	//				mul	$t0, $s4, $s3
memory[122] = 32'b00000001000010110100000000100001;	//				addu	$t0, $t0, $t3
memory[123] = 32'b00010110100000000000000000000100;	//				bne	$s4, $zero, irightnottop
memory[124] = 32'b00100110000010011111111111111111;	//				addiu	$t1, $s0, -1
memory[125] = 32'b01110001001100110100100000000010;	//				mul	$t1, $t1, $s3
memory[126] = 32'b00000001001010110100100000100001;	//				addu	$t1, $t1, $t3
memory[127] = 32'b00001000000000000000000010000111;	//				j	irightnotbottom
memory[128] = 32'b00100110100010011111111111111111;	//	irightnottop:		addiu	$t1, $s4, -1
memory[129] = 32'b01110001001100110100100000000010;	//				mul	$t1, $t1, $s3
memory[130] = 32'b00000001001010110100100000100001;	//				addu	$t1, $t1, $t3
memory[131] = 32'b00100110000010101111111111111111;	//	ifirightbottom:		addiu	$t2, $s0, -1
memory[132] = 32'b00010101010101000000000000000010;	//				bne	$t2, $s4, irightnotbottom
memory[133] = 32'b00000001011000000101000000100000;	//				add	$t2, $t3, $zero
memory[134] = 32'b00001000000000000000000010001010;	//				j	end
memory[135] = 32'b00100110100010100000000000000001;	//	irightnotbottom:	addiu	$t2, $s4, 1
memory[136] = 32'b01110001010100110101000000000010;	//				mul	$t2, $t2, $s3
memory[137] = 32'b00000001010010110101000000100001;	//				addu	$t2, $t2, $t3
memory[138] = 32'b00000000000010000100000010000000;	//	end:			sll	$t0, $t0, 2
memory[139] = 32'b00000000000010010100100010000000;	//				sll	$t1, $t1, 2
memory[140] = 32'b00000000000010100101000010000000;	//				sll	$t2, $t2, 2
memory[141] = 32'b00000001000001010100000000100001;	//				addu	$t0, $t0, $a1
memory[142] = 32'b00000001001001010100100000100001;	//				addu	$t1, $t1, $a1
memory[143] = 32'b00000001010001010101000000100001;	//				addu	$t2, $t2, $a1
memory[144] = 32'b10001101000011100000000000000000;	//				lw	$t6, 0($t0)
memory[145] = 32'b10001101001011010000000000000000;	//				lw	$t5, 0($t1)
memory[146] = 32'b10001101010011000000000000000000;	//				lw	$t4, 0($t2)
memory[147] = 32'b00010110101000000000000000010011;	//				bne	$s5, $zero, notleftcheckright
memory[148] = 32'b00110100000010000000000000000001;	//				ori	$t0, $zero, 1
memory[149] = 32'b00000001110010000111000000100100;	//				and	$t6, $t6, $t0
memory[150] = 32'b00000010111011101011100000100001;	//				addu	$s7, $s7, $t6
memory[151] = 32'b00000001101010000110100000100100;	//				and	$t5, $t5, $t0
memory[152] = 32'b00000010111011011011100000100001;	//				addu	$s7, $s7, $t5
memory[153] = 32'b00000001100010000110000000100100;	//				and	$t4, $t4, $t0
memory[154] = 32'b00000010111011001011100000100001;	//				addu	$s7, $s7, $t4
memory[155] = 32'b00111100000010001100000000000000;	//				lui	$t0, 49152
memory[156] = 32'b00000001111010000100100000100100;	//				and	$t1, $t7, $t0
memory[157] = 32'b00001100000000000000000100100101;	//				jal	countones
memory[158] = 32'b00000010111000101011100000100001;	//				addu	$s7, $s7, $v0
memory[159] = 32'b00000011000010000100100000100100;	//				and	$t1, $t8, $t0
memory[160] = 32'b00001100000000000000000100100101;	//				jal	countones
memory[161] = 32'b00000010111000101011100000100001;	//				addu	$s7, $s7, $v0
memory[162] = 32'b00111100000010000100000000000000;	//				lui	$t0, 16384
memory[163] = 32'b00000011001010000100100000100100;	//				and	$t1, $t9, $t0
memory[164] = 32'b00001100000000000000000100100101;	//				jal	countones
memory[165] = 32'b00000010111000101011100000100001;	//				addu	$s7, $s7, $v0
memory[166] = 32'b00001000000000000000000011001110;	//				j	markupdate
memory[167] = 32'b00110100000010000000000000011111;	//	notleftcheckright:	ori	$t0, $zero, 31
memory[168] = 32'b00010101000101010000000000010110;	//				bne	$t0, $s5, checkelse
memory[169] = 32'b00111100000010001000000000000000;	//				lui	$t0, 32768
memory[170] = 32'b00000001110010000100100000100100;	//				and	$t1, $t6, $t0
memory[171] = 32'b00001100000000000000000100100101;	//				jal	countones
memory[172] = 32'b00000010111000101011100000100001;	//				addu	$s7, $s7, $v0
memory[173] = 32'b00000001101010000100100000100100;	//				and	$t1, $t5, $t0
memory[174] = 32'b00001100000000000000000100100101;	//				jal	countones
memory[175] = 32'b00000010111000101011100000100001;	//				addu	$s7, $s7, $v0
memory[176] = 32'b00000001100010000100100000100100;	//				and	$t1, $t4, $t0
memory[177] = 32'b00001100000000000000000100100101;	//				jal	countones
memory[178] = 32'b00000010111000101011100000100001;	//				addu	$s7, $s7, $v0
memory[179] = 32'b00110100000010000000000000000011;	//				ori	$t0, $zero, 3
memory[180] = 32'b00000011000010000100100000100100;	//				and	$t1, $t8, $t0
memory[181] = 32'b00001100000000000000000100100101;	//				jal	countones
memory[182] = 32'b00000010111000101011100000100001;	//				addu	$s7, $s7, $v0
memory[183] = 32'b00000001111010000100100000100100;	//				and	$t1, $t7, $t0
memory[184] = 32'b00001100000000000000000100100101;	//				jal	countones
memory[185] = 32'b00000010111000101011100000100001;	//				addu	$s7, $s7, $v0
memory[186] = 32'b00110100000010000000000000000010;	//				ori	$t0, $zero, 2
memory[187] = 32'b00000011001010000100100000100100;	//				and	$t1, $t9, $t0
memory[188] = 32'b00001100000000000000000100100101;	//				jal	countones
memory[189] = 32'b00000010111000101011100000100001;	//				addu	$s7, $s7, $v0
memory[190] = 32'b00001000000000000000000011001110;	//				j	markupdate
memory[191] = 32'b00100010101010101111111111111111;	//	checkelse:		addi	$t2, $s5, -1
memory[192] = 32'b00111100000010001110000000000000;	//				lui	$t0, 57344
memory[193] = 32'b00000001010110000100100000000100;	//				sllv	$t1, $t8, $t2
memory[194] = 32'b00000001001010000100100000100100;	//				and	$t1, $t1, $t0
memory[195] = 32'b00001100000000000000000100100101;	//				jal	countones
memory[196] = 32'b00000010111000101011100000100001;	//				addu	$s7, $s7, $v0
memory[197] = 32'b00000001010011110100100000000100;	//				sllv	$t1, $t7, $t2
memory[198] = 32'b00000001001010000100100000100100;	//				and	$t1, $t1, $t0
memory[199] = 32'b00001100000000000000000100100101;	//				jal	countones
memory[200] = 32'b00000010111000101011100000100001;	//				addu	$s7, $s7, $v0
memory[201] = 32'b00111100000010001010000000000000;	//				lui	$t0, 40960
memory[202] = 32'b00000001010110010100100000000100;	//				sllv	$t1, $t9, $t2
memory[203] = 32'b00000001001010000100100000100100;	//				and	$t1, $t1, $t0
memory[204] = 32'b00001100000000000000000100100101;	//				jal	countones
memory[205] = 32'b00000010111000101011100000100001;	//				addu	$s7, $s7, $v0
memory[206] = 32'b00111100000010001000000000000000;	//	markupdate:		lui	$t0, 32768
memory[207] = 32'b00000010101010000100000000000110;	//				srlv	$t0, $t0, $s5
memory[208] = 32'b00000001000110010100000000100100;	//				and	$t0, $t0, $t9
memory[209] = 32'b00010101000000000000000000000110;	//				bne	$t0, $zero, notdead
memory[210] = 32'b00110100000010000000000000000011;	//				ori	$t0, $zero, 3
memory[211] = 32'b00010101000101110000000000000010;	//				bne	$t0, $s7, donotgrow
memory[212] = 32'b00110100000010110000000000000001;	//				ori	$t3, $zero, 1
memory[213] = 32'b00001000000000000000000011011111;	//				j	updatememory
memory[214] = 32'b00110100000010110000000000000000;	//	donotgrow:		ori	$t3, $zero, 0
memory[215] = 32'b00001000000000000000000011011111;	//				j	updatememory
memory[216] = 32'b00110100000010000000000000000010;	//	notdead:		ori	$t0, $zero, 2
memory[217] = 32'b00110100000010010000000000000011;	//				ori	$t1, $zero, 3
memory[218] = 32'b00010001000101110000000000000011;	//				beq	$t0, $s7, liveon
memory[219] = 32'b00010001001101110000000000000010;	//				beq	$t1, $s7, liveon
memory[220] = 32'b00110100000010110000000000000001;	//				ori	$t3, $zero, 1
memory[221] = 32'b00001000000000000000000011011111;	//				j	updatememory
memory[222] = 32'b00110100000010110000000000000000;	//	liveon:			ori	$t3, $zero, 0
memory[223] = 32'b01110010100100110100000000000010;	//	updatememory:		mul	$t0, $s4, $s3
memory[224] = 32'b00000001000101100100000000100001;	//				addu	$t0, $t0, $s6
memory[225] = 32'b00000000000010000100000010000000;	//				sll	$t0, $t0, 2
memory[226] = 32'b00000001000001100100000000100000;	//				add	$t0, $t0, $a2
memory[227] = 32'b10001101000010010000000000000000;	//				lw	$t1, 0($t0)
memory[228] = 32'b00000000000010010100100001000000;	//				sll	$t1, $t1, 1
memory[229] = 32'b00000001001010110100100000100000;	//				add	$t1, $t1, $t3
memory[230] = 32'b10101101000010010000000000000000;	//				sw	$t1, 0($t0)
memory[231] = 32'b00110100000101110000000000000000;	//				ori	$s7, $zero, 0
memory[232] = 32'b00110100000010000000000000100000;	//	nextbit:		ori	$t0, $zero, 32
memory[233] = 32'b00100110101101010000000000000001;	//				addiu	$s5, $s5, 1
memory[234] = 32'b00010101000101011111111100111000;	//				bne	$t0, $s5, getregisters
memory[235] = 32'b00110100000101010000000000000000;	//				ori	$s5, $zero, 0
memory[236] = 32'b00100110110101100000000000000001;	//				addiu	$s6, $s6, 1
memory[237] = 32'b00010110110100111111111100110000;	//				bne	$s6, $s3, getword
memory[238] = 32'b00110100000101100000000000000000;	//				ori	$s6, $zero, 0
memory[239] = 32'b00100110100101000000000000000001;	//				addiu	$s4, $s4, 1
memory[240] = 32'b00010110100100001111111100101101;	//				bne	$s4, $s0, getword
memory[241] = 32'b00110100000011010000000000000000;	//	updatelife:		ori	$t5, $zero, 0
memory[242] = 32'b01110010000100110111000000000010;	//				mul	$t6, $s0, $s3
memory[243] = 32'b00010001101011100000000000001001;	//	updatelifeloop:		beq	$t5, $t6, updatelifedone
memory[244] = 32'b00000000000011010100000010000000;	//				sll	$t0, $t5, 2
memory[245] = 32'b00000001000001010100100000100000;	//				add	$t1, $t0, $a1
memory[246] = 32'b00000001000001100101000000100000;	//				add	$t2, $t0, $a2
memory[247] = 32'b10001101001010110000000000000000;	//				lw	$t3, 0($t1)
memory[248] = 32'b10001101010011000000000000000000;	//				lw	$t4, 0($t2)
memory[249] = 32'b00000001100010110100000000100110;	//				xor	$t0, $t4, $t3
memory[250] = 32'b10101101001010000000000000000000;	//				sw	$t0, 0($t1)
memory[251] = 32'b00100001101011010000000000000001;	//				addi	$t5, $t5, 1
memory[252] = 32'b00001000000000000000000011110011;	//				j	updatelifeloop
memory[253] = 32'b00100110010100101111111111111111;	//	updatelifedone:		addiu	$s2, $s2, -1
memory[254] = 32'b00010110010000001111111100011011;	//				bne	$s2, $zero, generation
memory[255] = 32'b10001100100010000000000000001100;	//				lw	$t0, 12($a0)
memory[256] = 32'b10001100100110000000000000010000;	//				lw	$t8, 16($a0)
memory[257] = 32'b00100101000010101111111111111111;	//				addiu	$t2, $t0, -1
memory[258] = 32'b00110100000011100000000000000000;	//				ori	$t6, $zero, 0
memory[259] = 32'b01110001010100110101000000000010;	//				mul	$t2, $t2, $s3
memory[260] = 32'b00110100000011010000000000000000;	//				ori	$t5, $zero, 0
memory[261] = 32'b00000001010011100110000000100001;	//	countrowloop:		addu	$t4, $t2, $t6
memory[262] = 32'b00000000000011000110000010000000;	//				sll	$t4, $t4, 2
memory[263] = 32'b00000001100001010110000000100001;	//				addu	$t4, $t4, $a1
memory[264] = 32'b10001101100010010000000000000000;	//				lw	$t1, 0($t4)
memory[265] = 32'b00001100000000000000000100100101;	//				jal	countones
memory[266] = 32'b00000001101000100110100000100001;	//				addu	$t5, $t5, $v0
memory[267] = 32'b00100101110011100000000000000001;	//				addiu	$t6, $t6, 1
memory[268] = 32'b00010101110100111111111111111000;	//				bne	$t6, $s3, countrowloop
memory[269] = 32'b00000001101000000001000000100000;	//				add	$v0, $t5, $zero
memory[270] = 32'b00110100000010100000000000100000;	//				ori	$t2, $zero, 32
memory[271] = 32'b00110100000010111111111111111111;	//				ori	$t3, $zero, -1
memory[272] = 32'b00000011000000000110000000100000;	//				add	$t4, $t8, $zero
memory[273] = 32'b00000001100010100110000000100010;	//	locatecorrectcolumn:	sub	$t4, $t4, $t2
memory[274] = 32'b00100001011010110000000000000001;	//				addi	$t3, $t3, 1
memory[275] = 32'b00000000000011000000100000101010;	//				slt	$at, $zero, $t4
memory[276] = 32'b00010100001000001111111111111100;	//				bne	$at, $zero, locatecorrectcolumn
memory[277] = 32'b01110001010010110110000000000010;	//				mul	$t4, $t2, $t3
memory[278] = 32'b00000011000011001100000000100010;	//				sub	$t8, $t8, $t4
memory[279] = 32'b00000001010110001100000000100010;	//				sub	$t8, $t2, $t8
memory[280] = 32'b00110100000010000000000000000000;	//				ori	$t0, $zero, 0
memory[281] = 32'b00110100000110010000000000000001;	//				ori	$t9, $zero, 1
memory[282] = 32'b01110001000100110110000000000010;	//	countcolumnloop:	mul	$t4, $t0, $s3
memory[283] = 32'b00000001100010110110000000100001;	//				addu	$t4, $t4, $t3
memory[284] = 32'b00000000000011000110000010000000;	//				sll	$t4, $t4, 2
memory[285] = 32'b00000001100001010110000000100001;	//				addu	$t4, $t4, $a1
memory[286] = 32'b10001101100011000000000000000000;	//				lw	$t4, 0($t4)
memory[287] = 32'b00000011000011000110000000000110;	//				srlv	$t4, $t4, $t8
memory[288] = 32'b00000001100110010110000000100100;	//				and	$t4, $t4, $t9
memory[289] = 32'b00000000011011000001100000100000;	//				add	$v1, $v1, $t4
memory[290] = 32'b00100001000010000000000000000001;	//				addi	$t0, $t0, 1
memory[291] = 32'b00010101000100001111111111110110;	//				bne	$t0, $s0, countcolumnloop
memory[292] = 32'b00001000000000000000000100100100;	//	doneloop:		j	doneloop
memory[293] = 32'b00110100000000100000000000000000;	//	countones:		ori	$v0, $zero, 0
memory[294] = 32'b00010001001000000000000000000100;	//	countonesloop:		beq	$t1, $zero, countonesexit
memory[295] = 32'b00100101001010111111111111111111;	//				addiu	$t3, $t1, -1
memory[296] = 32'b00000001001010110100100000100100;	//				and	$t1, $t1, $t3
memory[297] = 32'b00100100010000100000000000000001;	//				addiu	$v0, $v0, 1
memory[298] = 32'b00001000000000000000000100100110;	//				j	countonesloop
memory[299] = 32'b00000011111000000000000000001000;	//	countonesexit:		jr	$ra

	
/*memory[0] = 32'b00000000000000000000000000000000;
memory[1] = 32'b00100011101111011111111111111100;	//	main:			addi	$sp, $sp, -4
memory[2] = 32'b10101111101111110000000000000000;	//				sw	$ra, 0($sp)
memory[3] = 32'b00110100000001000000000000000000;	//				ori	$a0, $zero, 0
memory[4] = 32'b00110100000001010000000000010100;	//				ori	$a1, $zero, 20
memory[5] = 32'b00001100000000000000000000001010;	//				jal	GOL
memory[6] = 32'b10001111101111110000000000000000;	//				lw	$ra, 0($sp)
memory[7] = 32'b00000000000000000000000000000000;	//				jr	$ra
memory[8] = 32'b00110100000111010000101011110000;	//	End:			nop
//memory[8] = 32'b00000000000000000000000000000000;	//				nop
memory[9] = 32'b00001000000000000000000000000111;	//				j	End
memory[10] = 32'b00110100000000100000000000000000;	//	GOL:			ori	$v0, $zero, 0
memory[11] = 32'b00110100000000110000000000000000;	//				ori	$v1, $zero, 0
memory[12] = 32'b00110100000010001111111011010100;	//				ori	$t0, $zero, -600
memory[13] = 32'b00000000000010000100000010000000;	//				sll	$t0, $t0, 2
memory[14] = 32'b00000011101010001110100000100000;	//				add	$sp, $sp, $t0
memory[15] = 32'b00000011101000000011000000100000;	//				add	$a2, $sp, $zero
memory[16] = 32'b00000011101010001110100000100000;	//				add	$sp, $sp, $t0
memory[17] = 32'b00000011101000000011100000100000;	//				add	$a3, $sp, $zero
memory[18] = 32'b10001100100100000000000000000000;	//				lw	$s0, 0($a0)
memory[19] = 32'b10001100100100010000000000000100;	//				lw	$s1, 4($a0)
memory[20] = 32'b10001100100100100000000000001000;	//				lw	$s2, 8($a0)
memory[21] = 32'b10001100100100110000000000001100;	//				lw	$s3, 12($a0)
memory[22] = 32'b10001100100101000000000000010000;	//				lw	$s4, 16($a0)
memory[23] = 32'b00100011101111011111111111110000;	//				addi	$sp, $sp, -16
memory[24] = 32'b10101111101111110000000000000000;	//				sw	$ra, 0($sp)
memory[25] = 32'b10101111101100100000000000000100;	//				sw	$s2, 4($sp)
memory[26] = 32'b10101111101100110000000000001000;	//				sw	$s3, 8($sp)
memory[27] = 32'b10101111101101000000000000001100;	//				sw	$s4, 12($sp)
memory[28] = 32'b00001100000000000000000000110001;	//				jal	CreateArray
memory[29] = 32'b10001111101111110000000000000000;	//				lw	$ra, 0($sp)
memory[30] = 32'b10001111101100100000000000000100;	//				lw	$s2, 4($sp)
memory[31] = 32'b10001111101100110000000000001000;	//				lw	$s3, 8($sp)
memory[32] = 32'b10001111101101000000000000001100;	//				lw	$s4, 12($sp)
memory[33] = 32'b00100011101111010000000000010000;	//				addi	$sp, $sp, 16
memory[34] = 32'b00100011101111011111111111111100;	//				addi	$sp, $sp, -4
memory[35] = 32'b10101111101111110000000000000000;	//				sw	$ra, 0($sp)
memory[36] = 32'b00001100000000000000000001010101;	//				jal	GenerationUpdate
memory[37] = 32'b10001111101111110000000000000000;	//				lw	$ra, 0($sp)
memory[38] = 32'b00100011101111010000000000000100;	//				addi	$sp, $sp, 4
memory[39] = 32'b00100011101111011111111111111100;	//				addi	$sp, $sp, -4
memory[40] = 32'b10101111101111110000000000000000;	//				sw	$ra, 0($sp)
memory[41] = 32'b00001100000000000000000011100101;	//				jal	CountLiving
memory[42] = 32'b10001111101111110000000000000000;	//				lw	$ra, 0($sp)
memory[43] = 32'b00100011101111010000000000000100;	//				addi	$sp, $sp, 4
memory[44] = 32'b00110100000010000000000000110011;	//				ori	$t0, $zero, 400
memory[45] = 32'b00000000000010000100000010000000;	//				sll	$t0, $t0, 2
memory[46] = 32'b00000011101010001110100000100000;	//				add	$sp, $sp, $t0
memory[47] = 32'b00000011101010001110100000100000;	//				add	$sp, $sp, $t0
memory[48] = 32'b00000011111000000000000000001000;	//				jr	$ra
memory[49] = 32'b00110100000010000000000000000000;	//	CreateArray:		ori	$t0, $zero, 0
memory[50] = 32'b00110100000010010000000000000000;	//				ori	$t1, $zero, 0
memory[51] = 32'b00110100000010100000000000000000;	//				ori	$t2, $zero, 0
memory[52] = 32'b00110100000010110000000000000000;	//				ori	$t3, $zero, 0
memory[53] = 32'b00100001000011000000000000000001;	//	CAOutFor:		addi	$t4, $t0, 1
memory[54] = 32'b00000000000100010110100101000010;	//				srl	$t5, $s1, 5
memory[55] = 32'b01110001100011010101000000000010;	//				mul	$t2, $t4, $t5
memory[56] = 32'b00110100000010010000000000000000;	//				ori	$t1, $zero, 0
memory[57] = 32'b01110001000100010110000000000010;	//	CAInFor:		mul	$t4, $t0, $s1
memory[58] = 32'b00000001100100010110000000100000;	//				add	$t4, $t4, $s1
memory[59] = 32'b00100001100011001111111111111111;	//				addi	$t4, $t4, -1
memory[60] = 32'b00000001100010011100000000100010;	//				sub	$t8, $t4, $t1
memory[61] = 32'b00000011000001110110100000100000;	//				add	$t5, $t8, $a3
memory[62] = 32'b10100001101000000000000000000000;	//				sb	$zero, 0($t5)
memory[63] = 32'b00000000000010010110000101000010;	//	CAIf1:			srl	$t4, $t1, 5
memory[64] = 32'b00110100000011010000000000100000;	//				ori	$t5, $zero, 32
memory[65] = 32'b01110001100011010110000000000010;	//				mul	$t4, $t4, $t5
memory[66] = 32'b00000001001011000110000000100010;	//				sub	$t4, $t1, $t4
memory[67] = 32'b00010101100000000000000000000100;	//				bne	$t4, $zero, CAIf2
memory[68] = 32'b00100001010010101111111111111111;	//				addi	$t2, $t2, -1
memory[69] = 32'b00000000000010100110000010000000;	//				sll	$t4, $t2, 2
memory[70] = 32'b00000001100001010110000000100000;	//				add	$t4, $t4, $a1
memory[71] = 32'b10001101100010110000000000000000;	//				lw	$t3, 0($t4)
memory[72] = 32'b00110100000011110000000000000001;	//	CAIf2:			ori	$t7, $zero, 1
memory[73] = 32'b00000001011011110110100000100100;	//				and	$t5, $t3, $t7
memory[74] = 32'b00000011000001100110000000100000;	//				add	$t4, $t8, $a2
memory[75] = 32'b00010101111011010000000000000010;	//				bne	$t7, $t5, CAElse
memory[76] = 32'b10100001100011110000000000000000;	//				sb	$t7, 0($t4)
memory[77] = 32'b00001000000000000000000001001111;	//				j	CAAfterElse
memory[78] = 32'b10100001100000000000000000000000;	//	CAElse:			sb	$zero, 0($t4)
memory[79] = 32'b00000000000010110101100001000010;	//	CAAfterElse:		srl	$t3, $t3, 1
memory[80] = 32'b00100001001010010000000000000001;	//				addi	$t1, $t1, 1
memory[81] = 32'b00010101001100011111111111100111;	//				bne	$t1, $s1, CAInFor///
memory[82] = 32'b00100001000010000000000000000001;	//				addi	$t0, $t0, 1
memory[83] = 32'b00010101000100001111111111100001;	//				bne	$t0, $s0, CAOutFor ///
memory[84] = 32'b00000011111000000000000000001000;	//				jr	$ra
memory[85] = 32'b00100011101111011111111111110000;	//	GenerationUpdate:	addi	$sp, $sp, -16
memory[86] = 32'b10101111101111110000000000000000;	//				sw	$ra, 0($sp)
memory[87] = 32'b10101111101100100000000000000100;	//				sw	$s2, 4($sp)
memory[88] = 32'b10101111101100110000000000001000;	//				sw	$s3, 8($sp)
memory[89] = 32'b10101111101101000000000000001100;	//				sw	$s4, 12($sp)
memory[90] = 32'b00001100000000000000000001101000;	//				jal	ScanArray
memory[91] = 32'b10001111101111110000000000000000;	//				lw	$ra, 0($sp)
memory[92] = 32'b10001111101100100000000000000100;	//				lw	$s2, 4($sp)
memory[93] = 32'b10001111101100110000000000001000;	//				lw	$s3, 8($sp)
memory[94] = 32'b10001111101101000000000000001100;	//				lw	$s4, 12($sp)
memory[95] = 32'b00100011101111010000000000010000;	//				addi	$sp, $sp, 16
memory[96] = 32'b00100011101111011111111111111100;	//				addi	$sp, $sp, -4
memory[97] = 32'b10101111101111110000000000000000;	//				sw	$ra, 0($sp)
memory[98] = 32'b00001100000000000000000011010110;	//				jal	UpdateArray
memory[99] = 32'b10001111101111110000000000000000;	//				lw	$ra, 0($sp)
memory[100] = 32'b00100011101111010000000000000100;	//				addi	$sp, $sp, 4
memory[101] = 32'b00100010010100101111111111111111;	//				addi	$s2, $s2, -1
memory[102] = 32'b00010110010000001111111111101110;	//				bne	$s2, $zero, GenerationUpdate///
memory[103] = 32'b00000011111000000000000000001000;	//				jr	$ra
memory[104] = 32'b00110100000100100000000000000000;	//	ScanArray:		ori	$s2, $zero, 0
memory[105] = 32'b00110100000100110000000000000000;	//				ori	$s3, $zero, 0
memory[106] = 32'b01110010000100011011000000000010;	//				mul	$s6, $s0, $s1
memory[107] = 32'b00110100000101110000000000000000;	//				ori	$s7, $zero, 0
memory[108] = 32'b00110100000101000000000000000000;	//				ori	$s4, $zero, 0
memory[109] = 32'b00000010010100010100000000100010;	//	SAFor:			sub	$t0, $s2, $s1
memory[110] = 32'b00100001000010001111111111111111;	//				addi	$t0, $t0, -1
memory[111] = 32'b00000010010100010100100000100010;	//				sub	$t1, $s2, $s1
memory[112] = 32'b00000010010100010101000000100010;	//				sub	$t2, $s2, $s1
memory[113] = 32'b00100001010010100000000000000001;	//				addi	$t2, $t2, 1
memory[114] = 32'b00100010010010111111111111111111;	//				addi	$t3, $s2, -1
memory[115] = 32'b00100010010011000000000000000001;	//				addi	$t4, $s2, 1
memory[116] = 32'b00000010010100010110100000100000;	//				add	$t5, $s2, $s1
memory[117] = 32'b00100001101011011111111111111111;	//				addi	$t5, $t5, -1
memory[118] = 32'b00000010010100010111000000100000;	//				add	$t6, $s2, $s1
memory[119] = 32'b00000010010100010111100000100000;	//				add	$t7, $s2, $s1
memory[120] = 32'b00100001111011110000000000000001;	//				addi	$t7, $t7, 1
memory[121] = 32'b00000010010100011100100000101010;	//	SAIf1:			slt	$t9, $s2, $s1
memory[122] = 32'b00010011001000000000000000000100;	//				beq	$t9, $zero, SAElseIf1
memory[123] = 32'b00000001000101100100000000100000;	//				add	$t0, $t0, $s6
memory[124] = 32'b00000001001101100100100000100000;	//				add	$t1, $t1, $s6
memory[125] = 32'b00000001010101100101000000100000;	//				add	$t2, $t2, $s6
memory[126] = 32'b00001000000000000000000010000110;	//				j	SAIf2
memory[127] = 32'b00100010000110001111111111111111;	//	SAElseIf1:		addi	$t8, $s0, -1
memory[128] = 32'b01110011000100011100000000000010;	//				mul	$t8, $t8, $s1
memory[129] = 32'b00000010010110001100000000101010;	//				slt	$t8, $s2, $t8
memory[130] = 32'b00010111000000000000000000000011;	//				bne	$t8, $zero, SAIf2
memory[131] = 32'b00000001101101100110100000100010;	//				sub	$t5, $t5, $s6
memory[132] = 32'b00000001110101100111000000100010;	//				sub	$t6, $t6, $s6
memory[133] = 32'b00000001111101100111100000100010;	//				sub	$t7, $t7, $s6
memory[134] = 32'b01110010111100011100000000000010;	//	SAIf2:			mul	$t8, $s7, $s1
memory[135] = 32'b00000010010110001100000000100010;	//				sub	$t8, $s2, $t8
memory[136] = 32'b00010111000000000000000000000011;	//				bne	$t8, $zero, SAIf3
memory[137] = 32'b00000001000100010100000000100000;	//				add	$t0, $t0, $s1
memory[138] = 32'b00000001011100010101100000100000;	//				add	$t3, $t3, $s1
memory[139] = 32'b00000001101100010110100000100000;	//				add	$t5, $t5, $s1
memory[140] = 32'b00100010111110000000000000000001;	//	SAIf3:			addi	$t8, $s7, 1
memory[141] = 32'b01110011000100011100000000000010;	//				mul	$t8, $t8, $s1
memory[142] = 32'b00000011000100101100000000100010;	//				sub	$t8, $t8, $s2
memory[143] = 32'b00110100000110010000000000000001;	//				ori	$t9, $zero, 1
memory[144] = 32'b00010111000110010000000000000011;	//				bne	$t8, $t9, SAIf4
memory[145] = 32'b00000001010100010101000000100010;	//				sub	$t2, $t2, $s1
memory[146] = 32'b00000001100100010110000000100010;	//				sub	$t4, $t4, $s1
memory[147] = 32'b00000001111100010111100000100010;	//				sub	$t7, $t7, $s1
memory[148] = 32'b00000001000001100100000000100000;	//	SAIf4:			add	$t0, $t0, $a2
memory[149] = 32'b00000001001001100100100000100000;	//				add	$t1, $t1, $a2
memory[150] = 32'b00000001010001100101000000100000;	//				add	$t2, $t2, $a2
memory[151] = 32'b00000001011001100101100000100000;	//				add	$t3, $t3, $a2
memory[152] = 32'b00000001100001100110000000100000;	//				add	$t4, $t4, $a2
memory[153] = 32'b00000001101001100110100000100000;	//				add	$t5, $t5, $a2
memory[154] = 32'b00000001110001100111000000100000;	//				add	$t6, $t6, $a2
memory[155] = 32'b00000001111001100111100000100000;	//				add	$t7, $t7, $a2
memory[156] = 32'b10000001000010000000000000000000;	//				lb	$t0, 0($t0)
memory[157] = 32'b10000001001010010000000000000000;	//				lb	$t1, 0($t1)
memory[158] = 32'b10000001010010100000000000000000;	//				lb	$t2, 0($t2)
memory[159] = 32'b10000001011010110000000000000000;	//				lb	$t3, 0($t3)
memory[160] = 32'b10000001100011000000000000000000;	//				lb	$t4, 0($t4)
memory[161] = 32'b10000001101011010000000000000000;	//				lb	$t5, 0($t5)
memory[162] = 32'b10000001110011100000000000000000;	//				lb	$t6, 0($t6)
memory[163] = 32'b10000001111011110000000000000000;	//				lb	$t7, 0($t7)
memory[164] = 32'b00000001000010011001100000100000;	//				add	$s3, $t0, $t1
memory[165] = 32'b00000010011010101001100000100000;	//				add	$s3, $s3, $t2
memory[166] = 32'b00000010011010111001100000100000;	//				add	$s3, $s3, $t3
memory[167] = 32'b00000010011011001001100000100000;	//				add	$s3, $s3, $t4
memory[168] = 32'b00000010011011011001100000100000;	//				add	$s3, $s3, $t5
memory[169] = 32'b00000010011011101001100000100000;	//				add	$s3, $s3, $t6
memory[170] = 32'b00000010011011111001100000100000;	//				add	$s3, $s3, $t7
memory[171] = 32'b00000010010001100100000000100000;	//				add	$t0, $s2, $a2
memory[172] = 32'b10000001000010000000000000000000;	//				lb	$t0, 0($t0)
memory[173] = 32'b00010000000010000000000000000010;	//				beq	$zero, $t0, SEQ1
memory[174] = 32'b00110100000010000000000000000000;	//				ori	$t0, $zero, 0
memory[175] = 32'b00010000000000000000000000000001;	//				beq	$zero, $zero, SEQ0
memory[176] = 32'b00110100000010000000000000000001;	//	SEQ1:			ori	$t0, $zero, 1
memory[177] = 32'b00110100000010010000000000000011;	//	SEQ0:			ori	$t1, $zero, 3
memory[178] = 32'b00010010011010010000000000000010;	//				beq	$s3, $t1, Seq1
memory[179] = 32'b00110100000010010000000000000000;	//				ori	$t1, $zero, 0
memory[180] = 32'b00010000000000000000000000000001;	//				beq	$zero, $zero, Seq0
memory[181] = 32'b00110100000010010000000000000001;	//	Seq1:			ori	$t1, $zero, 1
memory[182] = 32'b00000001000010010100000000100100;	//	Seq0:			and	$t0, $t0, $t1
memory[183] = 32'b00110100000010010000000000000001;	//				ori	$t1, $zero, 1
memory[184] = 32'b00010101001100110000000000000010;	//				bne	$t1, $s3, SLE1
memory[185] = 32'b00110100000010100000000000000001;	//				ori	$t2, $0, 1
memory[186] = 32'b00010000000000000000000000000001;	//				beq	$0, $0, SLE0
memory[187] = 32'b00000010011010010101000000101010;	//	SLE1:			slt	$t2, $s3, $t1
memory[188] = 32'b00110100000010010000000000000100;	//	SLE0:			ori	$t1, $zero, 4
memory[189] = 32'b00010101001100110000000000000010;	//				bne	$t1, $s3, SGE1
memory[190] = 32'b00110100000010110000000000000001;	//				ori	$t3, $0, 1
memory[191] = 32'b00010000000000000000000000000001;	//				beq	$0, $0, SGE0
memory[192] = 32'b00000001001100110101100000101010;	//	SGE1:			slt	$t3, $t1, $s3
memory[193] = 32'b00000001010010110100100000100101;	//	SGE0:			or	$t1, $t2, $t3
memory[194] = 32'b00000010010001100101000000100000;	//				add	$t2, $s2, $a2
memory[195] = 32'b10000001010010100000000000000000;	//				lb	$t2, 0($t2)
memory[196] = 32'b00110100000010110000000000000001;	//				ori	$t3, $zero, 1
memory[197] = 32'b00010001011010100000000000000010;	//				beq	$t3, $t2, SSeq1
memory[198] = 32'b00110100000010100000000000000000;	//				ori	$t2, $0, 0
memory[199] = 32'b00010000000000000000000000000001;	//				beq	$0, $0, SSeq0
memory[200] = 32'b00110100000010100000000000000001;	//	SSeq1:			ori	$t2, $0, 1
memory[201] = 32'b00000001001010100100100000100100;	//	SSeq0:			and	$t1, $t1, $t2
memory[202] = 32'b00000001000010010100000000100101;	//				or	$t0, $t0, $t1
memory[203] = 32'b00010001000000000000000000000011;	//				beq	$t0, $zero, SAEndLoop
memory[204] = 32'b00000010010001110100000000100000;	//				add	$t0, $s2, $a3
memory[205] = 32'b00110100000010010000000000000001;	//				ori	$t1, $zero, 1
memory[206] = 32'b10100001000010010000000000000000;	//				sb	$t1, 0($t0)
memory[207] = 32'b00100010010100100000000000000001;	//	SAEndLoop:		addi	$s2, $s2, 1
memory[208] = 32'b00100010100101000000000000000001;	//				addi	$s4, $s4, 1
memory[209] = 32'b00010110100100010000000000000010;	//				bne	$s4, $s1, Nots7increment
memory[210] = 32'b00100010111101110000000000000001;	//				addi	$s7, $s7, 1
memory[211] = 32'b00110100000101000000000000000000;	//				ori	$s4, $zero, 0
memory[212] = 32'b00010110010101101111111110011000;	//	Nots7increment:		bne	$s2, $s6, SAFor
memory[213] = 32'b00000011111000000000000000001000;	//				jr	$ra
memory[214] = 32'b00110100000010000000000000000000;	//	UpdateArray:		ori	$t0, $zero, 0
memory[215] = 32'b00110100000110000000000000000001;	//				ori	$t8, $zero, 1
memory[216] = 32'b00000001000001110100100000100000;	//	UAFor:			add	$t1, $t0, $a3
memory[217] = 32'b10000001001010010000000000000000;	//				lb	$t1, 0($t1)
memory[218] = 32'b00110100000010100000000000000001;	//				ori	$t2, $zero, 1
memory[219] = 32'b00010101001010100000000000000110;	//				bne	$t1, $t2, UAEndFor
memory[220] = 32'b00000001000001100100100000100000;	//				add	$t1, $t0, $a2
memory[221] = 32'b10000001001010100000000000000000;	//				lb	$t2, 0($t1)
memory[222] = 32'b00000001010110000101000000100110;	//				xor	$t2, $t2, $t8
memory[223] = 32'b10100001001010100000000000000000;	//				sb	$t2, 0($t1)
memory[224] = 32'b00000001000001110101000000100000;	//				add	$t2, $t0, $a3
memory[225] = 32'b10100001010000000000000000000000;	//				sb	$zero, 0($t2)
memory[226] = 32'b00100001000010000000000000000001;	//	UAEndFor:		addi	$t0, $t0, 1
memory[227] = 32'b00010101000101101111111111110100;	//				bne	$t0, $s6, UAFor ///
memory[228] = 32'b00000011111000000000000000001000;	//				jr	$ra
memory[229] = 32'b00110100000010000000000000000000;	//	CountLiving:		ori	$t0, $zero, 0
memory[230] = 32'b00100010011010011111111111111111;	//	CLFor1:			addi	$t1, $s3, -1
memory[231] = 32'b01110001001100010100100000000010;	//				mul	$t1, $t1, $s1
memory[232] = 32'b00000001001010000100100000100000;	//				add	$t1, $t1, $t0
memory[233] = 32'b00000001001001100100100000100000;	//				add	$t1, $t1, $a2
memory[234] = 32'b10000001001010010000000000000000;	//				lb	$t1, 0($t1)
memory[235] = 32'b00000000010010010001000000100000;	//				add	$v0, $v0, $t1
memory[236] = 32'b00100001000010000000000000000001;	//				addi	$t0, $t0, 1
memory[237] = 32'b00010101000100011111111111111000;	//				bne	$t0, $s1, CLFor1///
memory[238] = 32'b00110100000010000000000000000000;	//				ori	$t0, $zero, 0
memory[239] = 32'b00100010100010011111111111111111;	//	CLFor2:			addi	$t1, $s4, -1
memory[240] = 32'b01110001000100010101000000000010;	//				mul	$t2, $t0, $s1
memory[241] = 32'b00000001001010100100100000100000;	//				add	$t1, $t1, $t2
memory[242] = 32'b00000001001001100100100000100000;	//				add	$t1, $t1, $a2
memory[243] = 32'b10000001001010010000000000000000;	//				lb	$t1, 0($t1)
memory[244] = 32'b00000000011010010001100000100000;	//				add	$v1, $v1, $t1
memory[245] = 32'b00100001000010000000000000000001;	//				addi	$t0, $t0, 1
memory[246] = 32'b00010101000100001111111111111000;	//				bne	$t0, $s0, CLFor2///
memory[247] = 32'b00000011111000000000000000001000;	//				jr	$ra
*/

	end
	
	
	assign Instruction = memory[Address[31:2]];
	
	

endmodule
